
//------------------------------------------------------------------------------
// "rom.v"
//
// Authors : K. Nguyen 10/2015 (UCL)
//
//
//------------------------------------------------------------------------------
module rom (
	input	wire 		HCLK,
	input	wire		HRESETn,
	
	input  	wire [12:0]	addr,
	output 	wire [31:0]	rdata,
	input	wire 		cs
);
	//----------------------------------------------------------------------------------
	//	REG & WIRES :
	//----------------------------------------------------------------------------------
	reg [31:0] mem [0:8191];
  reg [31:0] mem_last;
	//----------------------------------------------------------------------------------
	//	ROM :
	//----------------------------------------------------------------------------------
	initial begin
		$readmemh("./../src/sw/code.hex", mem);
	end
	
  always @(posedge HCLK)
  begin
    mem_last <= cs  ? mem[addr] : 32'b0;
  end
	assign rdata = mem_last;//(cs & mem_sel) ? mem[addr] : 32'b0;
	
endmodule